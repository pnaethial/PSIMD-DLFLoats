`timescale 1ns/1ps

module PSIMD_tb;

    // Testbench Signals
    logic clk;
    logic rst_n;
    logic [31:0] instr;
    logic [63:0] rs1_core;
    logic [3:0] invalid;
    logic [3:0] inexact;
    logic [3:0] overflow;
    logic [3:0] underflow;
    logic [3:0] div_by_zero;
    logic [63:0] data_out_to_mem;
    logic [63:0] data_in_from_mem;
    logic [63:0] address;
    logic mem_read,mem_write;
    logic [63:0]data_out_1;
    logic [63:0]data1,data2,data3;

    PSIMD dut (
        .clk(clk),
        .rst_n(rst_n),
        .instr(instr),
        .rs1_core(rs1_core),
        .invalid(invalid),
        .inexact(inexact),
        .overflow(overflow),
        .underflow(underflow),
        .div_by_zero(div_by_zero),
        .data_out_to_mem(data_out_to_mem),
        .data1(data1),
        .data2(data2),
        .data3(data3),
        .data_in_from_mem(data_in_from_mem),
        .address(address),
        .mem_read(mem_read),
        .mem_write(mem_write),
        .data_out_1(data_out_1)
        );

    // Clock Generation
    always #25 clk = ~clk; // 10ns period clock

    // Test Procedure
    initial begin
        clk = 0;
        rst_n = 0;
        instr = 32'b000000000000_00000_000_00001_0001011;
        rs1_core = 32'b000000000000_00000_000_00000_0000000;
        
        #100;

        instr = 32'b000000001000_00000_000_00010_0001011;
        rs1_core = 32'b000000000000_00000_000_00000_0000000;
        
        #100;

        instr = 32'b000000010000_00000_000_00011_0001011;
        rs1_core = 32'b000000000000_00000_000_00000_0000000;

        #100;

        instr = 32'b000000011000_00000_000_00100_0001011;
        rs1_core = 32'b000000000000_00000_000_00000_0000000;
        #100;

        instr = 32'b000000101000_00000_000_00101_0001011;
        rs1_core = 32'b000000000000_00000_000_00000_0000000;
        #100;

        instr = 32'b000000110000_00000_000_00110_0001011;
        rs1_core = 32'b000000000000_00000_000_00000_0000000;
        
        #100;

        instr = 32'b000000111000_00000_000_00111_0001011;
        rs1_core = 32'b000000000000_00000_000_00000_0000000;
        
        #100;

        instr = 32'b000001000000_00000_000_01000_0001011;
        rs1_core = 32'b000000000000_00000_000_00000_0000000;
        
        #100;

        instr = 32'b000001001000_00000_000_01001_0001011;
        rs1_core = 32'b000000000000_00000_000_00000_0000000;
        
        #100;

        instr = 32'b000001010000_00000_000_01010_0001011;
        rs1_core = 32'b000000000000_00000_000_00000_0000000;
        
        #100;

        instr = 32'b000001011000_00000_000_01011_0001011;
        rs1_core = 32'b000000000000_00000_000_00000_0000000;
        
        #100;

        instr = 32'b000001100000_00000_000_01100_0001011;
        rs1_core = 32'b000000000000_00000_000_00000_0000000;
        
//       //store
//       #100;
//        instr = 32'b0000000_00000_00000_000_00000_0101011;
//        #100;
//        instr = 32'b0000000_00001_00000_000_01000_0101011;
//        #100;
//        instr = 32'b0000000_00010_00000_000_10000_0101011;
//        #100;
//        instr = 32'b0000000_00011_00000_000_11000_0101011;
//        #100;
//        instr = 32'b0000001_00100_00000_000_00000_0101011;
//        #100;
//        instr = 32'b0000001_00101_00000_000_01000_0101011;
//        #100;
//        instr = 32'b0000001_00110_00000_000_10000_0101011;
//        #100;
//        instr = 32'b0000001_00111_00000_000_11000_0101011;
//        #100;
//        instr = 32'b0000010_01000_00000_000_00000_0101011;
//        #100;
//        instr = 32'b0000010_01001_00000_000_01000_0101011;
//        #100
       
        
        //add       
       #100;
       instr = 32'b00000_00_00010_00001_000_00000_1011011;
       #100;
       instr = 32'b00000_00_00010_00001_000_00001_1011011;
       #100;
       instr = 32'b00000_00_00001_00011_000_00010_1011011;
       #100;
       instr = 32'b00000_00_00110_00101_000_00100_1011011;
       #100;
       instr = 32'b00000_00_00111_00100_000_00101_1011011;
       #100;
       instr = 32'b00000_00_00110_00111_000_00110_1011011;
       #100;
       instr = 32'b00000_00_01000_00000_000_00111_1011011;
       #100;
       instr = 32'b00000_00_01001_00010_000_01000_1011011;
       #100;
       instr = 32'b00000_00_00111_00001_000_01001_1011011;
       #100;
       instr = 32'b00000_00_01000_00001_000_01010_1011011;
//       #100;
//       instr = 32'b00000_00_00000_01000_011_01011_1011011;
//       #100;
//       instr = 32'b00000_00_00110_00101_001_01100_1011011;
//       #100;
//       instr = 32'b00000_00_00100_01001_010_01101_1011011;
//       #100;
//       instr = 32'b00000_00_00001_00101_000_01110_1011011;
       
       

//        //sub
//       #100;
//       instr = 32'b00001_00_00000_00001_000_00000_1011011;
//       #100;
//       instr = 32'b00001_00_00010_00001_001_00001_1011011;
//       #100;
//       instr = 32'b00001_00_00001_00011_010_00010_1011011;
//       #100;
//       instr = 32'b00001_00_00110_00101_100_00100_1011011;
//       #100;
//       instr = 32'b00001_00_00111_00100_101_00101_1011011;
//       #100;
//       instr = 32'b00001_00_00110_00111_110_00110_1011011;
//       #100;
//       instr = 32'b00001_00_01000_00000_111_00111_1011011;
//       #100;
//       instr = 32'b00001_00_01001_00010_011_01000_1011011;
//       #100;
//       instr = 32'b00001_00_00111_00001_010_01001_1011011;
//       #100;
//       instr = 32'b00001_00_01000_00001_101_01010_1011011;
//       #100;
//       instr = 32'b00001_00_00000_01000_011_01011_1011011;
//       #100;
//       instr = 32'b00001_00_00110_00101_000_01100_1011011;
//       #100;
//       instr = 32'b00001_00_00100_01001_001_01101_1011011;
//       #100;
//       instr = 32'b00001_00_00001_00101_000_01110_1011011;;

//      //mul
//       #100;
//       instr = 32'b00010_00_00000_00001_000_00000_1011011;
//       #100;
//       instr = 32'b00010_00_00010_00001_001_00001_1011011;
//       #100;
//       instr = 32'b00010_00_00001_00011_010_00010_1011011;
//       #100;
//       instr = 32'b00010_00_00110_00101_100_00100_1011011;
//       #100;
//       instr = 32'b00010_00_00111_00100_101_00101_1011011;
//       #100;
//       instr = 32'b00010_00_00110_00111_110_00110_1011011;
//       #100;
//       instr = 32'b00010_00_01000_00000_111_00111_1011011;
//       #100;
//       instr = 32'b00010_00_01001_00010_010_01000_1011011;
//       #100;
//       instr = 32'b00010_00_00111_00001_100_01001_1011011;
//       #100;
//       instr = 32'b00010_00_01000_00001_010_01010_1011011;
//       #100;
//       instr = 32'b00010_00_00000_01000_110_01011_1011011;
//       #100;
//       instr = 32'b00010_00_00110_00101_000_01100_1011011;
//       #100;
//       instr = 32'b00010_00_00100_01001_110_01101_1011011;
//       #100;
//       instr = 32'b00010_00_00001_00101_000_01110_1011011;
        
//        //div
//        #100;
//       instr = 32'b00011_00_00000_00001_000_00000_1011011;
//       #100;
//       instr = 32'b00011_00_00010_00001_001_00001_1011011;
//       #100;
//       instr = 32'b00011_00_00001_00011_010_00010_1011011;
//       #100;
//       instr = 32'b00011_00_00110_00101_011_00100_1011011;
//       #100;
//       instr = 32'b00011_00_00111_00100_100_00101_1011011;
//       #100;
//       instr = 32'b00011_00_00110_00111_101_00110_1011011;
//       #100;
//       instr = 32'b00011_00_01000_00000_110_00111_1011011;
//       #100;
//       instr = 32'b00011_00_01001_00010_111_01000_1011011;
//       #100;
//       instr = 32'b00011_00_00111_00001_101_01001_1011011;
//       #100;
//       instr = 32'b00011_00_01000_00001_110_01010_1011011;
//       #100;
//       instr = 32'b00011_00_00000_01000_001_01011_1011011;
//       #100;
//       instr = 32'b00011_00_00110_00101_010_01100_1011011;
//       #100;
//       instr = 32'b00011_00_00100_01001_110_01101_1011011;
//       #100;
//       instr = 32'b00011_00_00001_00101_010_01110_1011011;
        
        
//        #100;
//        instr = 32'b00011_00_00011_00001_000_00100_1011011;
        

//        //sqrt
//       #100;
//       instr = 32'b01011_00_00000_00001_000_00000_1011011;
//       #100;
//       instr = 32'b01011_00_00010_00001_001_00001_1011011;
//       #100;
//       instr = 32'b01011_00_00001_00011_010_00010_1011011;
//       #100;
//       instr = 32'b01011_00_00110_00101_011_00100_1011011;
//       #100;
//       instr = 32'b01011_00_00111_00100_100_00101_1011011;
//       #100;
//       instr = 32'b01011_00_00110_00111_101_00110_1011011;
//       #100;
//       instr = 32'b01011_00_01000_00000_110_00111_1011011;
//       #100;
//       instr = 32'b01011_00_01001_00010_111_01000_1011011;
//       #100;
//       instr = 32'b01011_00_00111_00001_001_01001_1011011;
//       #100;
//       instr = 32'b01011_00_01000_00001_010_01010_1011011;
//       #100;
//       instr = 32'b01011_00_00000_01000_110_01011_1011011;
//       #100;
//       instr = 32'b01011_00_00110_00101_010_01100_1011011;
//       #100;
//       instr = 32'b01011_00_00100_01001_011_01101_1011011;
//       #100;
//       instr = 32'b01011_00_00001_00101_010_01110_1011011;
        
//        //sign_inv
//       #100;
//       instr = 32'b00100_00_00000_00001_000_00000_1011011;
//       #100;
//       instr = 32'b000100_00_00010_00001_000_00001_1011011;
//       #100;
//       instr = 32'b00100_00_00001_00011_000_00010_1011011;
//       #100;
//       instr = 32'b00100_00_00110_00101_000_00100_1011011;
//       #100;
//       instr = 32'b00100_00_00111_00100_000_00101_1011011;
//       #100;
//       instr = 32'b00100_00_00110_00111_000_00110_1011011;
//       #100;
//       instr = 32'b00100_00_01000_00000_000_00111_1011011;
//       #100;
//       instr = 32'b00100_00_01001_00010_000_01000_1011011;
//       #100;
//       instr = 32'b00100_00_00111_00001_000_01001_1011011;
//       #100;
//       instr = 32'b00100_00_01000_00001_000_01010_1011011;
//       #100;
//       instr = 32'b00100_00_00000_01000_000_01011_1011011;
//       #100;
//       instr = 32'b00100_00_00110_00101_000_01100_1011011;
//       #100;
//       instr = 32'b00100_00_00100_01001_000_01101_1011011;
//       #100;
//       instr = 32'b00100_00_00001_00101_000_01110_1011011;
        
//        //sign_neg_inv
//      #100;
//       instr = 32'b00100_00_00000_00001_001_00000_1011011;
//       #100;
//       instr = 32'b00100_00_00010_00001_001_00001_1011011;
//       #100;
//       instr = 32'b00100_00_00001_00011_001_00010_1011011;
//       #100;
//       instr = 32'b00100_00_00110_00101_001_00100_1011011;
//       #100;
//       instr = 32'b00100_00_00111_00100_001_00101_1011011;
//       #100;
//       instr = 32'b00100_00_00110_00111_001_00110_1011011;
//       #100;
//       instr = 32'b00100_00_01000_00000_001_00111_1011011;
//       #100;
//       instr = 32'b00100_00_01001_00010_001_01000_1011011;
//       #100;
//       instr = 32'b00100_00_00111_00001_001_01001_1011011;
//       #100;
//       instr = 32'b00100_00_01000_00001_001_01010_1011011;
//       #100;
//       instr = 32'b00100_00_00000_01000_001_01011_1011011;
//       #100;
//       instr = 32'b00100_00_00110_00101_001_01100_1011011;
//       #100;
//       instr = 32'b00100_00_00100_01001_001_01101_1011011;
//       #100;
//       instr = 32'b00100_00_00001_00101_001_01110_1011011;
        
//        //sign xor
//       #100;
//       instr = 32'b00100_00_00000_00001_010_00000_1011011;
//       #100;
//       instr = 32'b00100_00_00010_00001_010_00001_1011011;
//       #100;
//       instr = 32'b00100_00_00001_00011_010_00010_1011011;
//       #100;
//       instr = 32'b00100_00_00110_00101_010_00100_1011011;
//       #100;
//       instr = 32'b00100_00_00111_00100_010_00101_1011011;
//       #100;
//       instr = 32'b00100_00_00110_00111_010_00110_1011011;
//       #100;
//       instr = 32'b00100_00_01000_00000_010_00111_1011011;
//       #100;
//       instr = 32'b00100_00_01001_00010_010_01000_1011011;
//       #100;
//       instr = 32'b00100_00_00111_00001_010_01001_1011011;
//       #100;
//       instr = 32'b00100_00_01000_00001_010_01010_1011011;
//       #100;
//       instr = 32'b00100_00_00000_01000_010_01011_1011011;
//       #100;
//       instr = 32'b00100_00_00110_00101_010_01100_1011011;
//       #100;
//       instr = 32'b00100_00_00100_01001_010_01101_1011011;
//       #100;
//       instr = 32'b00100_00_00001_00101_010_01110_1011011;
        
//        //min
//      #100;
//       instr = 32'b00101_00_00000_00001_000_00000_1011011;
//       #100;
//       instr = 32'b00101_00_00010_00001_000_00001_1011011;
//       #100;
//       instr = 32'b00101_00_00001_00011_000_00010_1011011;
//       #100;
//       instr = 32'b00101_00_00110_00101_000_00100_1011011;
//       #100;
//       instr = 32'b00101_00_00111_00100_000_00101_1011011;
//       #100;
//       instr = 32'b00101_00_00110_00111_000_00110_1011011;
//       #100;
//       instr = 32'b00101_00_01000_00000_000_00111_1011011;
//       #100;
//       instr = 32'b00101_00_01001_00010_000_01000_1011011;
//       #100;
//       instr = 32'b00101_00_00111_00001_000_01001_1011011;
//       #100;
//       instr = 32'b00101_00_01000_00001_000_01010_1011011;
//       #100;
//       instr = 32'b00101_00_00000_01000_000_01011_1011011;
//       #100;
//       instr = 32'b00101_00_00110_00101_000_01100_1011011;
//       #100;
//       instr = 32'b00101_00_00100_01001_000_01101_1011011;
//       #100;
//       instr = 32'b00101_00_00001_00101_000_01110_1011011;
        
//        //max
//      #100;
//       instr = 32'b00101_00_00000_00001_001_00000_1011011;
//       #100;
//       instr = 32'b00101_00_00010_00001_001_00001_1011011;
//       #100;
//       instr = 32'b00101_00_00001_00011_001_00010_1011011;
//       #100;
//       instr = 32'b00101_00_00110_00101_001_00100_1011011;
//       #100;
//       instr = 32'b00101_00_00111_00100_001_00101_1011011;
//       #100;
//       instr = 32'b00101_00_00110_00111_001_00110_1011011;
//       #100;
//       instr = 32'b00101_00_01000_00000_001_00111_1011011;
//       #100;
//       instr = 32'b00101_00_01001_00010_001_01000_1011011;
//       #100;
//       instr = 32'b00101_00_00111_00001_001_01001_1011011;
//       #100;
//       instr = 32'b00101_00_01000_00001_001_01010_1011011;
//       #100;
//       instr = 32'b00101_00_00000_01000_001_01011_1011011;
//       #100;
//       instr = 32'b00101_00_00110_00101_001_01100_1011011;
//       #100;
//       instr = 32'b00101_00_00100_01001_001_01101_1011011;
//       #100;
//       instr = 32'b00101_00_00001_00101_001_01110_1011011;
        
//        //dl to int
//        #100;
//        instr = 32'b01000_00_00000_00000_000_10000_1011011;
//        #100;
//        instr = 32'b01000_00_00000_00001_000_10001_1011011;
//        #100;
//        instr = 32'b01000_00_00000_00010_000_10010_1011011;
//        #100;
//        instr = 32'b01000_00_00000_00011_000_10011_1011011;
//        #100;
//        instr = 32'b01000_00_00000_00100_000_10100_1011011;
//        #100;
//        instr = 32'b01000_00_00000_00101_000_10101_1011011;
//        #100;
//        instr = 32'b01000_00_00000_00110_000_10110_1011011;
//        #100;
//        instr = 32'b01000_00_00000_00111_000_10111_1011011;
//        #100;
//        instr = 32'b01000_00_00000_01000_000_01100_1011011;
//        #100;
//        instr = 32'b01000_00_00000_01001_000_11001_1011011;
//        #100;
//        instr = 32'b01000_00_00000_01010_000_11010_1011011;
//        #100;
//        instr = 32'b01000_00_00000_01011_000_11100_1011011;
        
        
//        //int to dl
//       #100;
//        instr = 32'b01001_00_00000_00000_000_10000_1011011;
//        #100;
//        instr = 32'b01001_00_00000_00001_001_10001_1011011;
//        #100;
//        instr = 32'b01001_00_00000_00010_010_10010_1011011;
//        #100;
//        instr = 32'b01001_00_00000_00011_011_10011_1011011;
//        #100;
//        instr = 32'b01001_00_00000_00100_100_10100_1011011;
//        #100;
//        instr = 32'b01001_00_00000_00101_101_10101_1011011;
//        #100;
//        instr = 32'b01001_00_00000_00110_110_10110_1011011;
//        #100;
//        instr = 32'b01001_00_00000_00111_111_10111_1011011;
//        #100;
//        instr = 32'b01001_00_00000_01000_101_1100_1011011;
//        #100;
//        instr = 32'b01001_00_00000_01001_011_11001_1011011;
//        #100;
//        instr = 32'b01001_00_00000_01010_001_11010_1011011;
//        #100;
//        instr = 32'b01001_00_00000_01011_010_11100_1011011;
        
//        //equal
//      #100;
//       instr = 32'b10100_00_00000_00001_010_00000_1011011;
//       #100;
//       instr = 32'b10100_00_00010_00001_010_00001_1011011;
//       #100;
//       instr = 32'b10100_00_00001_00011_010_00010_1011011;
//       #100;
//       instr = 32'b10100_00_00110_00101_010_00100_1011011;
//       #100;
//       instr = 32'b10100_00_00111_00100_010_00101_1011011;
//       #100;
//       instr = 32'b10100_00_00110_00111_010_00110_1011011;
//       #100;
//       instr = 32'b10100_00_01000_00000_010_00111_1011011;
//       #100;
//       instr = 32'b10100_00_01001_00010_010_01000_1011011;
//       #100;
//       instr = 32'b10100_00_00111_00001_010_01001_1011011;
//       #100;
//       instr = 32'b10100_00_01000_00001_010_01010_1011011;
//       #100;
//       instr = 32'b10100_00_00000_01000_010_01011_1011011;
//       #100;
//       instr = 32'b10100_00_00110_00101_010_01100_1011011;
//       #100;
//       instr = 32'b10100_00_00100_01001_010_01101_1011011;
        
//        //less than
//      #100;
//       instr = 32'b10100_00_00000_00001_001_00000_1011011;
//       #100;
//       instr = 32'b10100_00_00010_00001_001_00001_1011011;
//       #100;
//       instr = 32'b10100_00_00001_00011_001_00010_1011011;
//       #100;
//       instr = 32'b10100_00_00110_00101_001_00100_1011011;
//       #100;
//       instr = 32'b10100_00_00111_00100_001_00101_1011011;
//       #100;
//       instr = 32'b10100_00_00110_00111_001_00110_1011011;
//       #100;
//       instr = 32'b10100_00_01000_00000_001_00111_1011011;
//       #100;
//       instr = 32'b10100_00_01001_00010_001_01000_1011011;
//       #100;
//       instr = 32'b10100_00_00111_00001_001_01001_1011011;
//       #100;
//       instr = 32'b10100_00_01000_00001_001_01010_1011011;
//       #100;
//       instr = 32'b10100_00_00000_01000_001_01011_1011011;
//       #100;
//       instr = 32'b10100_00_00110_00101_001_01100_1011011;
//       #100;
//       instr = 32'b10100_00_00100_01001_001_01101_1011011;
        
//        //less/equal
//       #100;
//       instr = 32'b10100_00_00000_00001_000_00000_1011011;
//       #100;
//       instr = 32'b10100_00_00010_00001_000_00001_1011011;
//       #100;
//       instr = 32'b10100_00_00001_00011_000_00010_1011011;
//       #100;
//       instr = 32'b10100_00_00110_00101_000_00100_1011011;
//       #100;
//       instr = 32'b10100_00_00111_00100_000_00101_1011011;
//       #100;
//       instr = 32'b10100_00_00110_00111_000_00110_1011011;
//       #100;
//       instr = 32'b10100_00_01000_00000_000_00111_1011011;
//       #100;
//       instr = 32'b10100_00_01001_00010_000_01000_1011011;
//       #100;
//       instr = 32'b10100_00_00111_00001_000_01001_1011011;
//       #100;
//       instr = 32'b10100_00_01000_00001_000_01010_1011011;
//       #100;
//       instr = 32'b10100_00_00000_01000_000_01011_1011011;
//       #100;
//       instr = 32'b10100_00_00110_00101_000_01100_1011011;
//       #100;
//       instr = 32'b10100_00_00100_01001_000_01101_1011011;
        
//        //mul add
//       #100;
//       instr = 32'b00000_00_00000_00001_000_00000_0011011;
//       #100;
//       instr = 32'b00010_00_00010_00001_000_00001_0011011;
//       #100;
//       instr = 32'b00001_00_00001_00011_001_00010_0011011;
//       #100;
//       instr = 32'b00011_00_00110_00101_010_00100_0011011;
//       #100;
//       instr = 32'b00100_00_00111_00100_100_00101_0011011;
//       #100;
//       instr = 32'b00101_00_00110_00111_011_00110_0011011;
//       #100;
//       instr = 32'b00110_00_01000_00000_101_00111_0011011;
//       #100;
//       instr = 32'b00111_00_01001_00010_110_01000_0011011;
//       #100;
//       instr = 32'b01000_00_00111_00001_111_01001_0011011;
//       #100;
//       instr = 32'b01001_00_01000_00001_010_01010_0011011;
//       #100;
//       instr = 32'b01010_00_00000_01000_110_01011_0011011;
//       #100;
//       instr = 32'b01011_00_00110_00101_011_01100_0011011;
//       #100;
//       instr = 32'b01100_00_00100_01001_001_01101_0011011;
//       #100;
//       instr = 32'b01101_00_00001_00101_101_01110_0011011;
        
//        //mul sub
//        #100;
//       instr = 32'b00000_00_00000_00001_000_00000_0111011;
//       #100;
//       instr = 32'b00010_00_00010_00001_000_00001_0111011;
//       #100;
//       instr = 32'b00001_00_00001_00011_001_00010_0111011;
//       #100;
//       instr = 32'b00011_00_00110_00101_010_00100_0111011;
//       #100;
//       instr = 32'b00100_00_00111_00100_100_00101_0111011;
//       #100;
//       instr = 32'b00101_00_00110_00111_111_00110_0111011;
//       #100;
//       instr = 32'b00110_00_01000_00000_110_00111_0111011;
//       #100;
//       instr = 32'b00111_00_01001_00010_010_01000_0111011;
//       #100;
//       instr = 32'b01000_00_00111_00001_011_01001_0111011;
//       #100;
//       instr = 32'b01001_00_01000_00001_100_01010_0111011;
//       #100;
//       instr = 32'b01010_00_00000_01000_110_01011_0111011;
//       #100;
//       instr = 32'b01011_00_00110_00101_011_01100_0111011;
//       #100;
//       instr = 32'b01100_00_00100_01001_001_01101_0111011;
//       #100;
//       instr = 32'b01101_00_00001_00101_000_01110_0111011;
        
       

        
        #100;
    $finish;
    end

endmodule
