`timescale 1ns / 1ps

module dlfloat16_decoder_tb;
  reg [31:0] instr;
  wire [3:0] ena;
  wire [2:0] rm;
  wire [2:0] sel2;
  wire op;
  wire [1:0] sel1;
  wire [4:0] rs1, rs2, rs3, rd;
  wire [11:0] imm;
  wire wr_enable;
  wire mem_read, mem_write, s_1, s_2,sp;

  dlfloat16_decoder uut (
    .instr(instr),
    .ena(ena),
    .rm(rm),
    .sel2(sel2),
    .op(op),
    .sel1(sel1),
    .rs1(rs1),
    .rs2(rs2),
    .rs3(rs3),
    .rd(rd),
    .imm(imm),
    .wr_enable(wr_enable),
    .mem_read(mem_read),
    .mem_write(mem_write),
    .s_1(s_1),
    .s_2(s_2),
    .sp(sp)
  );

  initial begin
//        //load
//        #10
//        instr = 32'b000000000000_00000_000_00000_0001011;
        
//        //store
//        #10
//        instr = 32'b0000000_01000_00000_000_00000_0101011;
        
        //add       
        #10
        instr = 32'b00000_00_00010_00001_000_00100_1011011;
        
       #100;
       instr = 32'b00000_00_00000_00001_000_00000_1011011;
       #100;
       instr = 32'b00000_00_00010_00001_001_00001_1011011;
       #100;
       instr = 32'b00000_00_00001_00011_010_00010_1011011;
       #100;
       instr = 32'b00000_00_00110_00101_011_00100_1011011;
       #100;
       instr = 32'b00000_00_00111_00100_100_00101_1011011;
       #100;
       instr = 32'b00000_00_00110_00111_101_00110_1011011;
       #100;
       instr = 32'b00000_00_01000_00000_110_00111_1011011;
        
//        //sub
//        #10
//        instr = 32'b00001_00_00011_00010_000_00100_1011011;
        
//        //mul
//        #10
//        instr = 32'b00010_00_00001_00000_000_00100_1011011;
        
//        //div
//        #10
//        instr = 32'b00011_00_00011_00010_000_00100_1011011;
        
//        //sqrt
//        #10
//        instr = 32'b01011_00_00000_00000_000_00100_1011011;
        
//        //sign_inv
//        #10
//        instr = 32'b00100_00_00011_00010_000_00100_1011011;
        
//        //sign_neg_inv
//        #10
//        instr = 32'b00100_00_00001_00000_001_00100_1011011;
        
//        //sign xor
//        #10
//        instr = 32'b00100_00_00011_00010_010_00100_1011011;
        
//        //min
//        #10
//        instr = 32'b00101_00_00001_00000_000_00100_1011011;
        
//        //max
//        #10
//        instr = 32'b00101_00_00011_00010_001_00100_1011011;
        
//        //dl to int
//        #10
//        instr = 32'b01000_00_00000_00000_000_00100_1011011;
        
//        //int to dl
//        #10
//        instr = 32'b01001_00_00000_00010_000_00100_1011011;
        
//        //equal
//        #10
//        instr = 32'b10100_00_00001_00000_010_00100_1011011;
        
//        //less than
//        #10
//        instr = 32'b10100_00_00011_00010_001_00100_1011011;
        
//        //less/equal
//        #10
//        instr = 32'b10100_00_00001_00000_000_00100_1011011;
        
//        //mul add
//        #10
//        instr = 32'b00100_00_00011_00010_000_00100_0011011;
        
//        //mul sub
//        #10
//        instr = 32'b00100_00_00001_00000_000_00100_0111011;
        
        #50
    
    $finish;
  end
endmodule
