module instr_buffer(
    input logic clk,
    output logic [31:0] instr
);

    logic [31:0] inst [35:0];
    logic i ;

initial begin
        inst[0] <= 32'b00000_00_00010_00001_000_00000_1011011;
        inst[1] <= 32'b00000_00_00010_00001_000_00001_1011011;
        inst[2] <= 32'b00001_00_00000_00001_000_00000_1011011;
        inst[3] <= 32'b00001_00_00001_00101_000_01110_1011011;
        inst[4] <= 32'b00010_00_00000_00001_000_00000_1011011;
        inst[5] <= 32'b00010_00_01000_00000_111_00111_1011011;
        inst[6] <= 32'b00011_00_00000_00001_000_00000_1011011;
        inst[7] <= 32'b00011_00_00110_00111_101_00110_1011011;
        inst[8] <= 32'b01011_00_00000_00001_000_00000_1011011;
        inst[9] <= 32'b01011_00_00111_00100_100_00101_1011011;
        inst[10] <= 32'b00100_00_00000_00001_000_00000_1011011;
        inst[11] <= 32'b00100_00_01000_00000_000_00111_1011011;
        inst[12] <= 32'b00100_00_00010_00001_001_00001_1011011;
        inst[13] <= 32'b00100_00_01000_00000_001_00111_1011011;
        inst[14] <= 32'b00100_00_00001_00011_010_00010_1011011;
        inst[15] <= 32'b00100_00_01000_00001_010_01010_1011011;
        inst[16] <= 32'b00101_00_00111_00001_000_01001_1011011;
        inst[17] <= 32'b00101_00_00110_00101_000_00100_1011011;
        inst[18] <= 32'b00101_00_00110_00101_001_00100_1011011;
        inst[19] <= 32'b00101_00_00111_00100_001_00101_1011011;
        inst[20] <= 32'b01000_00_00000_00101_000_10101_1011011;
        inst[21] <= 32'b01000_00_00000_01011_000_11100_1011011;
        inst[22] <= 32'b01001_00_00000_00001_001_10001_1011011;
        inst[23] <= 32'b01001_00_00000_01000_101_11000_1011011;
        inst[24] <= 32'b10100_00_01000_00000_010_00111_1011011;
        inst[25] <= 32'b10100_00_01000_00001_010_01010_1011011;
        inst[26] <= 32'b10100_00_00111_00100_001_00101_1011011;
        inst[27] <= 32'b10100_00_00000_01000_001_01011_1011011;
        inst[28] <= 32'b10100_00_00110_00111_000_00110_1011011;
        inst[29] <= 32'b10100_00_00111_00001_000_01001_1011011;
        inst[30] <= 32'b00100_00_00111_00100_100_00101_0011011;
        inst[31] <= 32'b00000_00_00000_00001_000_00000_0011011;
        inst[32] <= 32'b00100_00_00111_00100_100_00101_0111011;
        inst[33] <= 32'b01100_00_00100_01001_001_01101_0111011;
        
        i = 0;
end

always @(posedge clk) begin
        instr <= inst[i];
        if (i < 36)
            i <= i + 1;
end



endmodule
